// Listing 4.2
module d_ff_reset
   (
    input wire clk, reset,
    input wire d,
    output reg q
   );

   // body
   always @(posedge clk) begin
      if (reset) begin
         q <= 1'b0;
      end else begin
         q <= d;
      end
   end
endmodule
